package ibex_pkg_pext;

  //////////////////////
  // Multiplier modes //
  //////////////////////
  typedef enum logic[1:0] {
    M8x8, 
    M16x16, 
    M32x16, 
    M32x32
  } mult_pext_mode_e;

  ///////////////////////////
  // ALL P-ext instruxtion //
  ///////////////////////////
  typedef enum logic [7:0] {
    ZPN_ADD8,
    ZPN_ADD16,
    ZPN_ADD64,
    ZPN_AVE,
    ZPN_BITREV,
    ZPN_BITREVI,
    ZPN_BPICK,
    ZPN_CLROV,
    ZPN_CLRS8,
    ZPN_CLRS16,
    ZPN_CLRS32,
    ZPN_CLZ8,
    ZPN_CLZ16,
    ZPN_CLZ32,
    ZPN_CMPEQ8,
    ZPN_CMPEQ16,
    ZPN_CRAS16,
    ZPN_CRSA16,
    ZPN_INSB0,
    ZPN_INSB1,
    ZPN_INSB2,
    ZPN_INSB3,
    ZPN_KABS8,
    ZPN_KABS16,
    ZPN_KABSW,
    ZPN_KADD8,
    ZPN_KADD16,
    ZPN_KADD64,
    ZPN_KADDH,
    ZPN_KADDW,
    ZPN_KCRAS16,
    ZPN_KCRSA16,
    ZPN_KDMBB,
    ZPN_KDMBT,
    ZPN_KDMTT,
    ZPN_KDMABB,
    ZPN_KDMABT,
    ZPN_KDMATT,
    ZPN_KHM8,
    ZPN_KHMX8,
    ZPN_KHM16,
    ZPN_KHMX16,
    ZPN_KHMBB,
    ZPN_KHMBT,
    ZPN_KHMTT,
    ZPN_KMABB,
    ZPN_KMABT,
    ZPN_KMATT,
    ZPN_KMADA,
    ZPN_KMAXDA,
    ZPN_KMADS,
    ZPN_KMADRS,
    ZPN_KMAXDS,
    ZPN_KMAR64,
    ZPN_KMDA,
    ZPN_KMXDA,
    ZPN_KMMAC,
    ZPN_KMMACu,
    ZPN_KMMAWB,
    ZPN_KMMAWBu,
    ZPN_KMMAWB2,
    ZPN_KMMAWB2u,
    ZPN_KMMAWT,
    ZPN_KMMAWTu,
    ZPN_KMMAWT2,
    ZPN_KMMAWT2u,
    ZPN_KMMSB,
    ZPN_KMMSBu,
    ZPN_KMMWB2,
    ZPN_KMMWB2u,
    ZPN_KMMWT2,
    ZPN_KMMWT2u,
    ZPN_KMSDA,
    ZPN_KMSXDA,
    ZPN_KMSR64,
    ZPN_KSLLW,
    ZPN_KSLLIW,
    ZPN_KSLL8,
    ZPN_KSLLI8,
    ZPN_KSLL16,
    ZPN_KSLLI16,
    ZPN_KSLRA8,
    ZPN_KSLRA8u,
    ZPN_KSLRA16,
    ZPN_KSLRA16u,
    ZPN_KSLRAW,
    ZPN_KSLRAWu,
    ZPN_KSTAS16,
    ZPN_KSTSA16,
    ZPN_KSUB8,
    ZPN_KSUB16,
    ZPN_KSUB64,
    ZPN_KSUBH,
    ZPN_KSUBW,
    ZPN_KWMMUL,
    ZPN_KWMMULu,
    ZPN_MADDR32,
    ZPN_MAXW,
    ZPN_MINW,
    ZPN_MSUBR32,
    ZPN_MULR64,
    ZPN_MULSR64,
    ZPN_PBSAD,
    ZPN_PBSADA,
    ZPN_PKBB16,
    ZPN_PKBT16,
    ZPN_PKTT16,
    ZPN_PKTB16,
    ZPN_RADD8,
    ZPN_RADD16,
    ZPN_RADD64,
    ZPN_RADDW,
    ZPN_RCRAS16,
    ZPN_RCRSA16,
    ZPN_RDOV,
    ZPN_RSTAS16,
    ZPN_RSTSA16,
    ZPN_RSUB8,
    ZPN_RSUB16,
    ZPN_RSUB64,
    ZPN_RSUBW,
    ZPN_SCLIP8,
    ZPN_SCLIP16,
    ZPN_SCLIP32,
    ZPN_SCMPLE8,
    ZPN_SCMPLE16,
    ZPN_SCMPLT8,
    ZPN_SCMPLT16,
    ZPN_SLL8,
    ZPN_SLLI8,
    ZPN_SLL16,
    ZPN_SLLI16,
    ZPN_SMAL,
    ZPN_SMALBB,
    ZPN_SMALBT,
    ZPN_SMALTT,
    ZPN_SMALDA,
    ZPN_SMALXDA,
    ZPN_SMALDS,
    ZPN_SMALDRS,
    ZPN_SMALXDS,
    ZPN_SMAR64,
    ZPN_SMAQA,
    ZPN_SMAQAsu,
    ZPN_SMAX8,
    ZPN_SMAX16,
    ZPN_SMBB16,
    ZPN_SMBT16,
    ZPN_SMTT16,
    ZPN_SMDS,
    ZPN_SMDRS,
    ZPN_SMXDS,
    ZPN_SMIN8,
    ZPN_SMIN16,
    ZPN_SMMUL,
    ZPN_SMMULu,
    ZPN_SMMWB,
    ZPN_SMMWBu,
    ZPN_SMMWT,
    ZPN_SMMWTu,
    ZPN_SMSLDA,
    ZPN_SMSLXDA,
    ZPN_SMSR64,
    ZPN_SMUL8,
    ZPN_SMULX8,
    ZPN_SMUL16,
    ZPN_SMULX16,
    ZPN_SRAu,
    ZPN_SRAIu,
    ZPN_SRA8,
    ZPN_SRA8u,
    ZPN_SRAI8,
    ZPN_SRAI8u,
    ZPN_SRA16,
    ZPN_SRA16u,
    ZPN_SRAI16,
    ZPN_SRAI16u,
    ZPN_SRL8,
    ZPN_SRL8u,
    ZPN_SRLI8,
    ZPN_SRLI8u,
    ZPN_SRL16,
    ZPN_SRL16u,
    ZPN_SRLI16,
    ZPN_SRLI16u,
    ZPN_STAS16,
    ZPN_STSA16,
    ZPN_SUB8,
    ZPN_SUB16,
    ZPN_SUB64,
    ZPN_SUNPKD810,
    ZPN_SUNPKD820,
    ZPN_SUNPKD830,
    ZPN_SUNPKD831,
    ZPN_SUNPKD832,
    ZPN_SWAP8,
    ZPN_SWAP16,
    ZPN_UCLIP8,
    ZPN_UCLIP16,
    ZPN_UCLIP32,
    ZPN_UCMPLE8,
    ZPN_UCMPLE16,
    ZPN_UCMPLT8,
    ZPN_UCMPLT16,
    ZPN_UKADD8,
    ZPN_UKADD16,
    ZPN_UKADD64,
    ZPN_UKADDH,
    ZPN_UKADDW,
    ZPN_UKCRAS16,
    ZPN_UKCRSA16,
    ZPN_UKMAR64,
    ZPN_UKMSR64,
    ZPN_UKSTAS16,
    ZPN_UKSTSA16,
    ZPN_UKSUB8,
    ZPN_UKSUB16,
    ZPN_UKSUB64,
    ZPN_UKSUBH,
    ZPN_UKSUBW,
    ZPN_UMAR64,
    ZPN_UMAQA,
    ZPN_UMAX8,
    ZPN_UMAX16,
    ZPN_UMIN8,
    ZPN_UMIN16,
    ZPN_UMSR64,
    ZPN_UMUL8,
    ZPN_UMULX8,
    ZPN_UMUL16,
    ZPN_UMULX16,
    ZPN_URADD8,
    ZPN_URADD16,
    ZPN_URADD64,
    ZPN_URADDW,
    ZPN_URCRAS16,
    ZPN_URCRSA16,
    ZPN_URSTAS16,
    ZPN_URSTSA16,
    ZPN_URSUB8,
    ZPN_URSUB16,
    ZPN_URSUB64,
    ZPN_URSUBW,
    ZPN_WEXTI,
    ZPN_WEXT,
    ZPN_ZUNPKD810,
    ZPN_ZUNPKD820,
    ZPN_ZUNPKD830,
    ZPN_ZUNPKD831,
    ZPN_ZUNPKD832
  } zpn_op_e;

endpackage
